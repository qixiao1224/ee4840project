module vga_ball(input logic        clk,
	        input logic 	   reset,
		input logic [31:0]  writedata,
		input logic 	   write,
		input 		   chipselect,
		input logic [2:0]  address,

		output logic [7:0] VGA_R, VGA_G, VGA_B,
		output logic 	   VGA_CLK, VGA_HS, VGA_VS,
		                   VGA_BLANK_n,
		output logic 	   VGA_SYNC_n);

   logic [7:0] D0, D1, D2, D3, D4, C0, C1, C2, C3;
   logic [7:0] 	   background_r, background_g, background_b;
   logic [31:0] data_reg, control_reg;

   logic [10:0]	   hcount;
   logic [9:0]     vcount;

// vga_ball test
   logic [7:0] pos_v, pos_h;
   logic ball;
   logic [31:0] dish, disv;
   logic [10:0]   poshh;
   logic [9:0]    posvv;
   // One step is 16 bit
   assign poshh=pos_h<<4;
   assign posvv=pos_v<<4;
   // Calculate distance between current point and origin
   assign dish= (poshh[10:1] > hcount)?(poshh[10:1] - hcount[10:1]): (hcount[10:1] -poshh[10:1]); // hcount[10:1] is pixel column
   assign disv= (posvv > vcount)?(posvv - vcount): (vcount - posvv);
   assign ball = dish*dish+disv*disv < 16'd16 *16'd16;

// vga counter
   vga_counters counters(.clk50(clk), .*);

//wire between modules
logic [7:0] read_image0,read_image1,read_image2,read_image3,read_conv,read_dense;
logic [14:0] conv_ram_addr_a,conv_ram_addr_b,dense_ram_addr_a,dense_ram_addr_b;
logic [9:0] image_ram_addr_a,image_ram_addr_b;
logic we_image0,we_image1,we_image2,we_image3,we_conv,we_dense;
logic [7:0] data_image0,data_image1,data_image2,data_image3,data_conv,data_dense;

memory memory1( 
    .clk(clk),
    .reset(reset),

//input from image_ram
    //memory_read
    .image_ram_addr_b(image_ram_addr_b),
    //memory_write
    .image_ram_addr_a(image_ram_addr_a),
    .data_image0(data_image0),
    .data_image1(data_image1),
    .data_image2(data_image2),
    .data_image3(data_image3),
    .we_image0(we_image0),
    .we_image1(we_image1),
    .we_iamge2(we_image2),
    .we_image3(we_image3),

//input from conv_Ram
//memory_read
    .conv_ram_addr_b(conv_ram_addr_b),
//memory_write
    .conv_ram_addr_a(conv_ram_addr_a),
    .data_conv(data_conv),
    .we_conv(we_conv),

//input from dense_ram
//memory_read
.dense_ram_addr_b(conv_ram_addr_b),
//memory_write
    .dense_ram_addr_a(dense_ram_addr_a),
    .data_dense(data_dense),
    .we_dense(we_dense),

//outputs from RAM
//memory_read 
    .read_image0(read_image0), 
    .read_image1(read_image1), 
    .read_image2(read_image2), 
    .read_image3(read_image3),
    .read_conv(read_conv)
    .read_dense(read_dense),
);

memory_write memory_write1(
    .clk(clk),
    .reset(reset),
    .writedata(//TODO),
    .control_reg(//TODO),
    
    .wren0(we_image0),
    .wren1(we_image1),
    .wren2(we_image2),
    .wren3(we_image3),
    .wren_conv(we_conv),
    .wren_dense(we_conv),
    .data0(data_image0),
    .data1(data_image1),
    .data2(data_image2),
    .data3(data_image3),
    .data4(data_conv),
    .data5(data_dense),
    .image_ram_addr(image_ram_addr_a),
    .conv_ram_addr(conv_ram_addr_a),
    .dense_ram_addr(dense_ram_addr_a)
);



memory_read memory_read1(
    .clk(clk),
    .reset(reset),

    //read from outter ram
    .read_image0(read_image0), 
    .read_image1(read_image1), 
    .read_image2(read_image2), 
    .read_image3(read_image3),
    .read_conv(read_conv)
    .read_dense(read_dense),

    //TODO: NOT WIRED
    .out0(//TODO), 
    .out1(//TODO), 
    .out2(//TODO), 
    .out3(//TODO), 
    .out_param(//TODO),
    //output logic [7:0] filter0,filter1,filter2,filter3,

    //output read address to upper level
    .image_ram_addr(image_ram_addr_b);
    .conv_ram_addr(conv_ram_addr_b);
    .dense_ram_addr(dense_ram_addr_b);

);


   always_ff @(posedge clk)
     if (reset) begin
	background_r <= 8'h0;
	background_g <= 8'h0;
	background_b <= 8'h80;
	control_reg <= 0;
	data_reg <= 0;
	// vga_ball test
	pos_v <= 8'h0;
	pos_h <= 8'h0;
     end else if (chipselect && write) begin
		case (address)
			3'h0: begin
				control_reg <= writedata;
				data_reg <= 0;
				pos_v <= writedata[7:0];
				end
			3'h1: begin
				data_reg <= writedata;
				control_reg <= 0; // TODO Need to check
				pos_h <= writedata[7:0];
				end
		endcase
	end

   always_comb begin
      {VGA_R, VGA_G, VGA_B} = {8'h0, 8'h0, 8'h0};
      if (VGA_BLANK_n )
        if (ball) begin
	  {VGA_R, VGA_G, VGA_B} = {8'hff, 8'hff, 8'hff};
        end
	else
	  {VGA_R, VGA_G, VGA_B} =
             {background_r, background_g, background_b};
   end
	       

endmodule

module vga_counters(
 input logic 	     clk50, reset,
 output logic [10:0] hcount,  // hcount[10:1] is pixel column
 output logic [9:0]  vcount,  // vcount[9:0] is pixel row
 output logic 	     VGA_CLK, VGA_HS, VGA_VS, VGA_BLANK_n, VGA_SYNC_n);

/*
 * 640 X 480 VGA timing for a 50 MHz clock: one pixel every other cycle
 * 
 * HCOUNT 1599 0             1279       1599 0
 *             _______________              ________
 * ___________|    Video      |____________|  Video
 * 
 * 
 * |SYNC| BP |<-- HACTIVE -->|FP|SYNC| BP |<-- HACTIVE
 *       _______________________      _____________
 * |____|       VGA_HS          |____|
 */
   // Parameters for hcount
   parameter HACTIVE      = 11'd 1280,
             HFRONT_PORCH = 11'd 32,
             HSYNC        = 11'd 192,
             HBACK_PORCH  = 11'd 96,   
             HTOTAL       = HACTIVE + HFRONT_PORCH + HSYNC +
                            HBACK_PORCH; // 1600
   
   // Parameters for vcount
   parameter VACTIVE      = 10'd 480,
             VFRONT_PORCH = 10'd 10,
             VSYNC        = 10'd 2,
             VBACK_PORCH  = 10'd 33,
             VTOTAL       = VACTIVE + VFRONT_PORCH + VSYNC +
                            VBACK_PORCH; // 525

   logic endOfLine;
   
   always_ff @(posedge clk50 or posedge reset)
     if (reset)          hcount <= 0;
     else if (endOfLine) hcount <= 0;
     else  	         hcount <= hcount + 11'd 1;

   assign endOfLine = hcount == HTOTAL - 1;
       
   logic endOfField;
   
   always_ff @(posedge clk50 or posedge reset)
     if (reset)          vcount <= 0;
     else if (endOfLine)
       if (endOfField)   vcount <= 0;
       else              vcount <= vcount + 10'd 1;

   assign endOfField = vcount == VTOTAL - 1;

   // Horizontal sync: from 0x520 to 0x5DF (0x57F)
   // 101 0010 0000 to 101 1101 1111
   assign VGA_HS = !( (hcount[10:8] == 3'b101) &
		      !(hcount[7:5] == 3'b111));
   assign VGA_VS = !( vcount[9:1] == (VACTIVE + VFRONT_PORCH) / 2);

   assign VGA_SYNC_n = 1'b0; // For putting sync on the green signal; unused
   
   // Horizontal active: 0 to 1279     Vertical active: 0 to 479
   // 101 0000 0000  1280	       01 1110 0000  480
   // 110 0011 1111  1599	       10 0000 1100  524
   assign VGA_BLANK_n = !( hcount[10] & (hcount[9] | hcount[8]) ) &
			!( vcount[9] | (vcount[8:5] == 4'b1111) );

   /* VGA_CLK is 25 MHz
    *             __    __    __
    * clk50    __|  |__|  |__|
    *        
    *             _____       __
    * hcount[0]__|     |_____|
    */
   assign VGA_CLK = hcount[0]; // 25 MHz clock: rising edge sensitive
   
endmodule
